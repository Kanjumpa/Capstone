-- TX module that sends DATA when START is 1
-- BUSY: flag to show trasmission in progress


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


ENTITY TX IS
PORT(
	CLK: 	IN STD_LOGIC;
	START:		IN STD_LOGIC;
	BUSY:			OUT STD_LOGIC;
	DATA:			IN STD_LOGIC_VECTOR(17 downto 0);
	TX_LINE:		OUT STD_LOGIC
);
END TX;

ARCHITECTURE MAIN OF TX IS
SIGNAL PRSCL: INTEGER RANGE 0 TO 41667:=0;
SIGNAL INDEX: INTEGER RANGE 0 TO 30:=0;
SIGNAL DATAFLL: STD_LOGIC_VECTOR(17 downto 0);
SIGNAL TX_FLG: STD_LOGIC:='0';
BEGIN

PROCESS(CLK)
BEGIN
IF(CLK'EVENT AND CLK='1')THEN
	IF(TX_FLG='0' AND START='1')THEN
		TX_FLG<='1';
		BUSY<='1';
		DATAFLL <= DATA;
	END IF;
	
	IF(TX_FLG='1')THEN
		IF(PRSCL<5207)THEN
			PRSCL<=PRSCL+1;
		ELSE
			PRSCL<=0;
		END IF;
		
		IF(PRSCL=2604)THEN
			IF(INDEX=0)THEN
				TX_LINE<='1';
				INDEX<=1;
			ELSIF(INDEX=1)THEN
				TX_LINE<=DATAFLL(0);
				INDEX<=2;
			ELSIF(INDEX=2)THEN
				TX_LINE<=DATAFLL(1);
				INDEX<=3;
			ELSIF(INDEX=3)THEN
				TX_LINE<=DATAFLL(2);
				INDEX<=4;
			ELSIF(INDEX=4)THEN
				TX_LINE<=DATAFLL(3);
				INDEX<=5;
			ELSIF(INDEX=5)THEN
				TX_LINE<=DATAFLL(4);
				INDEX<=6;
			ELSIF(INDEX=6)THEN
				TX_LINE<=DATAFLL(5);
				INDEX<=7;
			ELSIF(INDEX=7)THEN
				TX_LINE<=DATAFLL(6);
				INDEX<=8;
			ELSIF(INDEX=8)THEN
				TX_LINE<=DATAFLL(7);
				INDEX<=9;
			ELSIF(INDEX=9)THEN
				TX_LINE<='1';
				INDEX<=10;
			ELSIF(INDEX=10)THEN
				TX_LINE<='0';
				INDEX<=11;
			ELSIF(INDEX=11)THEN
				TX_LINE<=DATAFLL(8);
				INDEX<=12;
			ELSIF(INDEX=12)THEN
				TX_LINE<=DATAFLL(9);
				INDEX<=13;
			ELSIF(INDEX=13)THEN
				TX_LINE<=DATAFLL(10);
				INDEX<=14;
			ELSIF(INDEX=14)THEN
				TX_LINE<=DATAFLL(11);
				INDEX<=15;
			ELSIF(INDEX=15)THEN
				TX_LINE<=DATAFLL(12);
				INDEX<=16;
			ELSIF(INDEX=16)THEN
				TX_LINE<=DATAFLL(13);
				INDEX<=17;
			ELSIF(INDEX=17)THEN
				TX_LINE<=DATAFLL(14);
				INDEX<=18;
			ELSIF(INDEX=18)THEN
				TX_LINE<=DATAFLL(15);
				INDEX<=19;
			ELSIF(INDEX=19)THEN
				TX_LINE<='1'; -- stop bit
				INDEX<=20;
			ELSIF(INDEX=20)THEN
				TX_LINE<='0'; -- start bit
				INDEX<=21;
			ELSIF(INDEX=21)THEN
				TX_LINE<=DATAFLL(16);
				INDEX<=22;
			ELSIF(INDEX=22)THEN
				TX_LINE<=DATAFLL(17);
				INDEX<=23;
			ELSIF(INDEX=23)THEN
				TX_LINE<='0';
				INDEX<=24;
			ELSIF(INDEX=24)THEN
				TX_LINE<='0';
				INDEX<=25;
			ELSIF(INDEX=25)THEN
				TX_LINE<='0';
				INDEX<=26;
			ELSIF(INDEX=26)THEN
				TX_LINE<='0';
				INDEX<=27;
			ELSIF(INDEX=27)THEN
				TX_LINE<='0';
				INDEX<=28;
			ELSIF(INDEX=28)THEN
				TX_LINE<='0';
				INDEX<=29;
			ELSIF(INDEX=29)THEN
				TX_LINE<='1'; -- stop bit
				INDEX<=30;
			ELSE
				TX_FLG<='0';
				BUSY<='0';
				INDEX<=0;
			END IF;	
		END IF;
	END IF;
END IF;
END PROCESS;
END MAIN;